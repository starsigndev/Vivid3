module Vivid.Test

class TestClass 

    func TestClass() 

        List ant;

        ant.Add(25);
        ant.Add(35);
        ant.Add(45.5);
        ant.Add(30.20);

        int a;

        foreach(a in ant)

            debug(a);

        end 

    end 

end 


