module Vivid.Test


class TestClass

  

    func TestClass()

        int a=0;

        for(a=0;a<50;a=a+1)

            debug(a);

        end 

    end 

end 


