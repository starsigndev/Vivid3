module Vivid.Test


class TestClass

    static int test=25;

    static func Other(int a)

        debug(a);

    end 

    func TestClass()

        TestClass.test = 85;

        TestClass.Other(20);



    end 

end 


