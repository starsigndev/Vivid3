module Vivid.Test

class CheckClass

end 

class TestClass

    int ant = 25;

    func TestClass()

        ant = 255*100;

        debug(ant);    

    end 

end 


