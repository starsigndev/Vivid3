module Vivid.Test


class TestClass

  
    func TestClass() 

      float a = 7;

       for(a=0;a<100;a=a+0.1)

            debug(a); : a<40;

        end 

    end 

end 


