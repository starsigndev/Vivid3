module Vivid.Maths.Vec3

class Vec3

    float X,Y,Z;

    func Vec3()

        X=0.0;
        Y=0.0;
        Z=0.0;

    end 

end 

