module Vivid.Game

class GameScript

    Node node;

    func GameScript()

        node = new Node();
        Debug("Game Script!");

    end 

  

end     