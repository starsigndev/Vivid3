module Vivid.Maths.Vec3

class Vec4

    CObj C;

    func Vec4()

        

    end 

end 

