module Vivid.Test

class TestClass

    int ant,other,cool;

    func TestClass(int my,int other,int test)

    end 

end 


