module Vivid.Test

class CheckClass

    int antony = 45;

    func CheckClass(int a)

       

    end 

end 

class TestClass


    func TestClass()

        CheckClass ant = new CheckClass(5);
        
        ant.antony = 100;

        debug(ant.antony+30); 

    end 

end 


