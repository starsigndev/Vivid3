module Vivid.Maths.Matrix4

class Matrix

    CObject C;

    func Matrix()

    end 

end 