module Vivid.Test

class TestClass

    int check = 1200,other;

    func test(int a)

       debug(a);

    end

    func TestClass()

        test(255);

    end 

end 


